module sort;
    reg power, clk, load_word;
    reg [15:0] in_word;
    reg [15:0] in_address;

    subleq uut(.power(power), .clk(clk), .load_word(load_word), .in_word(in_word), .in_address(in_address));

    initial begin
        power = 0;
        clk = 0;
        load_word = 0;

        
        #10

        load_word = 1;

        #2
in_address = 16'b0000000000000001;
in_word = 16'b0000000100000000;
#2
in_address = 16'b0000000000000010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000000011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000000100;
in_word = 16'b0000000100001100;
#2
in_address = 16'b0000000000000101;
in_word = 16'b0000000100001100;
#2
in_address = 16'b0000000000000110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000000111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000001000;
in_word = 16'b0000000100001100;
#2
in_address = 16'b0000000000001001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000001010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000001011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000001100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000001101;
in_word = 16'b0000000100001011;
#2
in_address = 16'b0000000000001110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000001111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000010000;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000000010001;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000000010010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000010011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000010100;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000000010101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000010110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000010111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000011000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000011001;
in_word = 16'b0000000100000000;
#2
in_address = 16'b0000000000011010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000011011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000011100;
in_word = 16'b0000000100001101;
#2
in_address = 16'b0000000000011101;
in_word = 16'b0000000100001101;
#2
in_address = 16'b0000000000011110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000011111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000100000;
in_word = 16'b0000000100001101;
#2
in_address = 16'b0000000000100001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000100010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000100011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000100100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000100101;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000000100110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000100111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000101000;
in_word = 16'b0000000011000001;
#2
in_address = 16'b0000000000101001;
in_word = 16'b0000000011000001;
#2
in_address = 16'b0000000000101010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000101011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000101100;
in_word = 16'b0000000011000001;
#2
in_address = 16'b0000000000101101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000101110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000101111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000110000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000110001;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000000110010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000110011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000110100;
in_word = 16'b0000000011001101;
#2
in_address = 16'b0000000000110101;
in_word = 16'b0000000011001101;
#2
in_address = 16'b0000000000110110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000110111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000111000;
in_word = 16'b0000000011001101;
#2
in_address = 16'b0000000000111001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000111010;
in_word = 16'b0000000100001110;
#2
in_address = 16'b0000000000111011;
in_word = 16'b0000000011001101;
#2
in_address = 16'b0000000000111100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000111101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000111110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000000111111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001000000;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000001000001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001000010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001000011;
in_word = 16'b0000000011010000;
#2
in_address = 16'b0000000001000100;
in_word = 16'b0000000011010000;
#2
in_address = 16'b0000000001000101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001000110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001000111;
in_word = 16'b0000000011010000;
#2
in_address = 16'b0000000001001000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001001001;
in_word = 16'b0000000100001110;
#2
in_address = 16'b0000000001001010;
in_word = 16'b0000000011010000;
#2
in_address = 16'b0000000001001011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001001100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001001101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001001110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001001111;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000001010000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001010001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001010010;
in_word = 16'b0000000011010001;
#2
in_address = 16'b0000000001010011;
in_word = 16'b0000000011010001;
#2
in_address = 16'b0000000001010100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001010101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001010110;
in_word = 16'b0000000011010001;
#2
in_address = 16'b0000000001010111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001011000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001011001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001011010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001011011;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000001011100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001011101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001011110;
in_word = 16'b0000000011010011;
#2
in_address = 16'b0000000001011111;
in_word = 16'b0000000011010011;
#2
in_address = 16'b0000000001100000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001100001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001100010;
in_word = 16'b0000000011010011;
#2
in_address = 16'b0000000001100011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001100100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001100101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001100110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001100111;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000001101000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001101001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001101010;
in_word = 16'b0000000011010111;
#2
in_address = 16'b0000000001101011;
in_word = 16'b0000000011010111;
#2
in_address = 16'b0000000001101100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001101101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001101110;
in_word = 16'b0000000011010111;
#2
in_address = 16'b0000000001101111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001110000;
in_word = 16'b0000000100001110;
#2
in_address = 16'b0000000001110001;
in_word = 16'b0000000011010111;
#2
in_address = 16'b0000000001110010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001110011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001110100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001110101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001110110;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000001110111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001111000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001111001;
in_word = 16'b0000000011011001;
#2
in_address = 16'b0000000001111010;
in_word = 16'b0000000011011001;
#2
in_address = 16'b0000000001111011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001111100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001111101;
in_word = 16'b0000000011011001;
#2
in_address = 16'b0000000001111110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000001111111;
in_word = 16'b0000000100001110;
#2
in_address = 16'b0000000010000000;
in_word = 16'b0000000011011001;
#2
in_address = 16'b0000000010000001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010000010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010000011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010000100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010000101;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000010000110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010000111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010001000;
in_word = 16'b0000000011011010;
#2
in_address = 16'b0000000010001001;
in_word = 16'b0000000011011010;
#2
in_address = 16'b0000000010001010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010001011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010001100;
in_word = 16'b0000000011011010;
#2
in_address = 16'b0000000010001101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010001110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010001111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010010000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010010001;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000010010010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010010011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010010100;
in_word = 16'b0000000011011111;
#2
in_address = 16'b0000000010010101;
in_word = 16'b0000000011011111;
#2
in_address = 16'b0000000010010110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010010111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010011000;
in_word = 16'b0000000011011111;
#2
in_address = 16'b0000000010011001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010011010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010011011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010011100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010011101;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000010011110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010011111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010100000;
in_word = 16'b0000000011101000;
#2
in_address = 16'b0000000010100001;
in_word = 16'b0000000011101000;
#2
in_address = 16'b0000000010100010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010100011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010100100;
in_word = 16'b0000000011101000;
#2
in_address = 16'b0000000010100101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010100110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010100111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010101000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010101001;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000010101010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010101011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010101100;
in_word = 16'b0000000011101001;
#2
in_address = 16'b0000000010101101;
in_word = 16'b0000000011101001;
#2
in_address = 16'b0000000010101110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010101111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010110000;
in_word = 16'b0000000011101001;
#2
in_address = 16'b0000000010110001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010110010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010110011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010110100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010110101;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000010110110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010110111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010111000;
in_word = 16'b0000000011101100;
#2
in_address = 16'b0000000010111001;
in_word = 16'b0000000011101100;
#2
in_address = 16'b0000000010111010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010111011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010111100;
in_word = 16'b0000000011101100;
#2
in_address = 16'b0000000010111101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010111110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000010111111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011000000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011000001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011000010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011000011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011000100;
in_word = 16'b0000000011111101;
#2
in_address = 16'b0000000011000101;
in_word = 16'b0000000011111101;
#2
in_address = 16'b0000000011000110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011000111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011001000;
in_word = 16'b0000000011111101;
#2
in_address = 16'b0000000011001001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011001010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011001011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011001100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011001101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011001110;
in_word = 16'b0000000011111101;
#2
in_address = 16'b0000000011001111;
in_word = 16'b0000000011110001;
#2
in_address = 16'b0000000011010000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011010001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011010010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011010011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011010100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011010101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011010110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011010111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011011000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011011001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011011010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011011011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011011100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011011101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011011110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011011111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011100000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011100001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011100010;
in_word = 16'b0000000011111101;
#2
in_address = 16'b0000000011100011;
in_word = 16'b0000000011111101;
#2
in_address = 16'b0000000011100100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011100101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011100110;
in_word = 16'b0000000011111101;
#2
in_address = 16'b0000000011100111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011101000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011101001;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011101010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011101011;
in_word = 16'b0000000011111101;
#2
in_address = 16'b0000000011101100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011101101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011101110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011101111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011110000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011110001;
in_word = 16'b0000000100001110;
#2
in_address = 16'b0000000011110010;
in_word = 16'b0000000011111110;
#2
in_address = 16'b0000000011110011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011110100;
in_word = 16'b0000000100001110;
#2
in_address = 16'b0000000011110101;
in_word = 16'b0000000100001101;
#2
in_address = 16'b0000000011110110;
in_word = 16'b0000000000100101;
#2
in_address = 16'b0000000011110111;
in_word = 16'b0000000100001110;
#2
in_address = 16'b0000000011111000;
in_word = 16'b0000000100001100;
#2
in_address = 16'b0000000011111001;
in_word = 16'b0000000000001101;
#2
in_address = 16'b0000000011111010;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011111011;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011111100;
in_word = 16'b0000000011111010;

#2
in_address = 16'b0000000000000000;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011111101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011111110;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000011111111;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000100000000;
in_word = 16'b1111111111110111;
#2
in_address = 16'b0000000100000001;
in_word = 16'b0000000000001001;
#2
in_address = 16'b0000000100000010;
in_word = 16'b0000000000000011;
#2
in_address = 16'b0000000100000011;
in_word = 16'b0000000000000100;
#2
in_address = 16'b0000000100000100;
in_word = 16'b0000000000000001;
#2
in_address = 16'b0000000100000101;
in_word = 16'b0000000000010111;
#2
in_address = 16'b0000000100000110;
in_word = 16'b0000000000000101;
#2
in_address = 16'b0000000100000111;
in_word = 16'b0000000000000110;
#2
in_address = 16'b0000000100001000;
in_word = 16'b0000000000010011;
#2
in_address = 16'b0000000100001001;
in_word = 16'b0000000000000010;
#2
in_address = 16'b0000000100001010;
in_word = 16'b0000000000001010;
#2
in_address = 16'b0000000100001011;
in_word = 16'b0000000100000001;
#2
in_address = 16'b0000000100001100;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000100001101;
in_word = 16'b0000000000000000;
#2
in_address = 16'b0000000100001110;
in_word = 16'b1111111111111111;


        #10

        load_word = 0;

        power = 1;

        #1500
        $stop;
    end

    always #5 clk = ~clk;

endmodule
