`timescale 1ns / 1ps

module FourBitAdder(
	 input a4,
    input a3,
    input a2,
    input a1,
    input a0,
	 input b4,
    input b3,
    input b2,
    input b1,
    input b0,
    input carryIn,
    output s3,
    output s2,
    output s1,
    output s0,
    output carryOut
    );

wire b0prime;
wire 
FullAdder fa1();
wire 
FullAdder fa1();

endmodule
